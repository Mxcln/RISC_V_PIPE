
`include "define.v"

module  hazard(
    input   wire                arst_n  ,

    input   wire    ex_
);





    assign  hazard_hold_o = id_ex_mem_r_i & id_ex_

endmodule
